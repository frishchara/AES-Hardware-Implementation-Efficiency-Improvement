module GFM(a,b,c);

input [7:0] a,b;
output [7:0] c;

wire [7:0] w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13;

assign w0={8{a[7]}}&b;
assign w1={w0[6],w0[5],w0[4],w0[3],w0[2],w0[1],w0[0],1'b0}^{{8{w0[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w2=w1^{8{a[6]}}&b;
assign w3={w2[6],w2[5],w2[4],w2[3],w2[2],w2[1],w2[0],1'b0}^{{8{w2[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w4=w3^{8{a[5]}}&b;
assign w5={w4[6],w4[5],w4[4],w4[3],w4[2],w4[1],w4[0],1'b0}^{{8{w4[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w6=w5^{8{a[4]}}&b;
assign w7={w6[6],w6[5],w6[4],w6[3],w6[2],w6[1],w6[0],1'b0}^{{8{w6[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w8=w7^{8{a[3]}}&b;
assign w9={w8[6],w8[5],w8[4],w8[3],w8[2],w8[1],w8[0],1'b0}^{{8{w8[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w10=w9^{8{a[2]}}&b;
assign w11={w10[6],w10[5],w10[4],w10[3],w10[2],w10[1],w10[0],1'b0}^{{8{w10[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w12=w11^{8{a[1]}}&b;
assign w13={w12[6],w12[5],w12[4],w12[3],w12[2],w12[1],w12[0],1'b0}^{{8{w12[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign c=w13^{8{a[0]}}&b;

endmodule
