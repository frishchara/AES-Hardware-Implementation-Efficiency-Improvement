module SBox (
    input [7:0] B,
    output [7:0] D
);

    wire [7:0] M [7:0];
    assign M[0] = 8'b10001111;
    assign M[1] = 8'b11000111;
    assign M[2] = 8'b11100011;
    assign M[3] = 8'b11110001;
    assign M[4] = 8'b11111000;
    assign M[5] = 8'b01111100;
    assign M[6] = 8'b00111110;
    assign M[7] = 8'b00011111;
	 wire [7:0] b;     
	 
    wire [7:0] C[0:7];
    assign C[0] = 8'h1; assign C[1] = 8'h1; assign C[2] = 8'h0; assign C[3] = 8'h0;
    assign C[4] = 8'h0; assign C[5] = 8'h1; assign C[6] = 8'h1; assign C[7] = 8'h0;
	 
	 ninv n0(.I(B), .O(b));


    assign D[0] = (M[0][7] & b[0])^(M[0][6] & b[1])^(M[0][5] & b[2])^(M[0][4] & b[3])^(M[0][3] & b[4])^(M[0][2] & b[5])^(M[0][1] & b[6])^(M[0][0] & b[7]) ^ C[0];
    assign D[1] = (M[1][7] & b[0])^(M[1][6] & b[1])^(M[1][5] & b[2])^(M[1][4] & b[3])^(M[1][3] & b[4])^(M[1][2] & b[5])^(M[1][1] & b[6])^(M[1][0] & b[7]) ^ C[1];
    assign D[2] = (M[2][7] & b[0])^(M[2][6] & b[1])^(M[2][5] & b[2])^(M[2][4] & b[3])^(M[2][3] & b[4])^(M[2][2] & b[5])^(M[2][1] & b[6])^(M[2][0] & b[7]) ^ C[2];
    assign D[3] = (M[3][7] & b[0])^(M[3][6] & b[1])^(M[3][5] & b[2])^(M[3][4] & b[3])^(M[3][3] & b[4])^(M[3][2] & b[5])^(M[3][1] & b[6])^(M[3][0] & b[7]) ^ C[3];
    assign D[4] = (M[4][7] & b[0])^(M[4][6] & b[1])^(M[4][5] & b[2])^(M[4][4] & b[3])^(M[4][3] & b[4])^(M[4][2] & b[5])^(M[4][1] & b[6])^(M[4][0] & b[7]) ^ C[4];
    assign D[5] = (M[5][7] & b[0])^(M[5][6] & b[1])^(M[5][5] & b[2])^(M[5][4] & b[3])^(M[5][3] & b[4])^(M[5][2] & b[5])^(M[5][1] & b[6])^(M[5][0] & b[7]) ^ C[5];
    assign D[6] = (M[6][7] & b[0])^(M[6][6] & b[1])^(M[6][5] & b[2])^(M[6][4] & b[3])^(M[6][3] & b[4])^(M[6][2] & b[5])^(M[6][1] & b[6])^(M[6][0] & b[7]) ^ C[6];
    assign D[7] = (M[7][7] & b[0])^(M[7][6] & b[1])^(M[7][5] & b[2])^(M[7][4] & b[3])^(M[7][3] & b[4])^(M[7][2] & b[5])^(M[7][1] & b[6])^(M[7][0] & b[7]) ^ C[7];

endmodule
